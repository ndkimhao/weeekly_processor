-- ##############################################################
-- ## BEGIN UOPS ROM
-- ##############################################################

type TArrUopROM is array (0 to 200-1) of std_logic_vector(1+UopLen-1 downto 0);
constant uops_rom : TArrUopROM := (
	/*   0 */ 14x"0000", --     nop # dummy instruction at index 0 & 1
	/*   1 */ 14x"0000", --     nop, !FALLTHROUGH
	/*     */            -- # ======================================
	/*     */            -- # pre-boot code
	/*     */            -- reset:
	/*     */            --     # --------------------
	/*     */            --     # reset arch registers
	/*   2 */ 14x"0110", --     mov A,  0
	/*   3 */ 14x"0120", --     mov B,  0
	/*   4 */ 14x"0130", --     mov C,  0
	/*   5 */ 14x"0140", --     mov D,  0
	/*   6 */ 14x"0150", --     mov SP, 0
	/*   7 */ 14x"0160", --     mov PC, 0
	/*   8 */ 14x"0170", --     mov FL, 0
	/*     */            --     # --------------------
	/*     */            --     # reset MMU
	/*     */            --     # phy=A:B, idx=X, start=Y, end=Z
	/*   9 */ 14x"02b0", --     con K, 1
	/*  10 */ 14x"018b", --     mov X, K
	/*  11 */ 14x"0190", --     mov Y, 0
	/*  12 */ 14x"02a1", --     con Z, 0xFFFF
	/*  13 */ 14x"0300", --     mmu # idx=1, 0000-FFFF to 0000-FFFF
	/*  14 */ 14x"0291", --     con Y, 0xFFFF
	/*  15 */ 14x"01a0", --     mov Z, 0
	/*  16 */ 14x"0c8b", --     alu X, K, ADD
	/*  17 */ 14x"0300", --     mmu # idx=1
	/*  18 */ 14x"0212", --     con A, 0xFF # and B = 0
	/*  19 */ 14x"0293", --     con Y, 0xD000
	/*  20 */ 14x"02a1", --     con Z, 0xFFFF
	/*  21 */ 14x"0c8b", --     alu X, K, ADD
	/*  22 */ 14x"0300", --     mmu # idx=2
	/*  23 */ 14x"0110", --     mov A, 0
	/*  24 */ 14x"0291", --     con Y, 0xFFFF
	/*  25 */ 14x"01a0", --     mov Z, 0
	/*  26 */ 14x"0c8b", --     alu X, K, ADD
	/*  27 */ 14x"0300", --     mmu # idx=3
	/*  28 */ 14x"0000", --     nop # wait 1 cycle to write MMU config
	/*     */            --     # --------------------
	/*     */            --     # reset Fetcher
	/*  29 */ 14x"0160", --     mov PC, 0
	/*  30 */ 14x"2263", --     con PC, 0xD000
	/*     */            -- # ======================================
	/*     */            -- # ALU
	/*     */            -- alu_2dd:
	/*  31 */ 14x"0988", --     (2d-) arg X, GET_0
	/*  32 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  33 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  34 */ 14x"2888", --     (2d-) arg X, PUT
	/*     */            -- alu_2di:
	/*  35 */ 14x"0988", --     (2d-) arg X, GET_0
	/*  36 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  37 */ 14x"0499", --     (--i) mem Y, Y, LOAD
	/*  38 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  39 */ 14x"2888", --     (2d-) arg X, PUT
	/*     */            -- alu_2id:
	/*  40 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  41 */ 14x"048b", --     (2i-) mem X, K, LOAD
	/*  42 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  43 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  44 */ 14x"25b8", --     (2i-) mem K, X, STORE
	/*     */            -- alu_2ii:
	/*  45 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  46 */ 14x"048b", --     (2i-) mem X, K, LOAD
	/*  47 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  48 */ 14x"0499", --     (--i) mem Y, Y, LOAD
	/*  49 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  50 */ 14x"25b8", --     (2i-) mem K, X, STORE
	/*     */            -- alu_3dd:
	/*  51 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  52 */ 14x"0baa", --     (3--) arg Z, GET_2
	/*  53 */ 14x"0f9a", --     (3--) alu Y, Z, OP_COPY
	/*  54 */ 14x"2899", --     (3d-) arg Y, PUT
	/*     */            -- alu_3di:
	/*  55 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  56 */ 14x"0499", --     (--i) mem Y, Y, LOAD
	/*  57 */ 14x"0baa", --     (3--) arg Z, GET_2
	/*  58 */ 14x"0f9a", --     (3--) alu Y, Z, OP_COPY
	/*  59 */ 14x"2899", --     (3d-) arg Y, PUT
	/*     */            -- alu_3id:
	/*  60 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  61 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  62 */ 14x"0baa", --     (3--) arg Z, GET_2
	/*  63 */ 14x"0f9a", --     (3--) alu Y, Z, OP_COPY
	/*  64 */ 14x"25b9", --     (3i-) mem K, Y, STORE
	/*     */            -- alu_3ii:
	/*  65 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  66 */ 14x"0a99", --     (---) arg Y, GET_1
	/*  67 */ 14x"0499", --     (--i) mem Y, Y, LOAD
	/*  68 */ 14x"0baa", --     (3--) arg Z, GET_2
	/*  69 */ 14x"0f9a", --     (3--) alu Y, Z, OP_COPY
	/*  70 */ 14x"25b9", --     (3i-) mem K, Y, STORE
	/*     */            -- alu_single_1dx:
	/*  71 */ 14x"0988", --     (1d-) arg X, GET_0
	/*  72 */ 14x"0f88", --     (1--) alu X, X, OP_COPY
	/*  73 */ 14x"2888", --     (-d-) arg X, PUT
	/*     */            -- alu_single_1ix:
	/*  74 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  75 */ 14x"048b", --     (1i-) mem X, K, LOAD
	/*  76 */ 14x"0f88", --     (1--) alu X, X, OP_COPY
	/*  77 */ 14x"25b8", --     (-i-) mem K, X, STORE
	/*     */            -- alu_single_2dd:
	/*  78 */ 14x"0a99", --     (2--) arg Y, GET_1
	/*  79 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  80 */ 14x"2888", --     (-d-) arg X, PUT
	/*     */            -- alu_single_2di:
	/*  81 */ 14x"0a99", --     (2--) arg Y, GET_1
	/*  82 */ 14x"0499", --     (2-i) mem Y, Y, LOAD
	/*  83 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  84 */ 14x"2888", --     (-d-) arg X, PUT
	/*     */            -- alu_single_2id:
	/*  85 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  86 */ 14x"0a99", --     (2--) arg Y, GET_1
	/*  87 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  88 */ 14x"25b8", --     (-i-) mem K, X, STORE
	/*     */            -- alu_single_2ii:
	/*  89 */ 14x"09bb", --     (-i-) arg K, GET_0
	/*  90 */ 14x"0a99", --     (2--) arg Y, GET_1
	/*  91 */ 14x"0499", --     (2-i) mem Y, Y, LOAD
	/*  92 */ 14x"0f89", --     (2--) alu X, Y, OP_COPY
	/*  93 */ 14x"25b8", --     (-i-) mem K, X, STORE
	/*     */            -- # ======================================
	/*     */            -- # CMP
	/*     */            -- cmp_dd:
	/*  94 */ 14x"0988", --     (--) arg X, GET_0
	/*  95 */ 14x"0a99", --     (--) arg Y, GET_1
	/*  96 */ 14x"3289", --     (--) cmp X, Y, OP_COPY
	/*     */            -- cmp_di:
	/*  97 */ 14x"0988", --     (--) arg X, GET_0
	/*  98 */ 14x"0a99", --     (--) arg Y, GET_1
	/*  99 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 100 */ 14x"3289", --     (--) cmp X, Y, OP_COPY
	/*     */            -- cmp_id:
	/* 101 */ 14x"0988", --     (--) arg X, GET_0
	/* 102 */ 14x"0488", --     (i-) mem X, X, LOAD
	/* 103 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 104 */ 14x"3289", --     (--) cmp X, Y, OP_COPY
	/*     */            -- cmp_ii:
	/* 105 */ 14x"0988", --     (--) arg X, GET_0
	/* 106 */ 14x"0488", --     (i-) mem X, X, LOAD
	/* 107 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 108 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 109 */ 14x"3289", --     (--) cmp X, Y, OP_COPY
	/*     */            -- # ======================================
	/*     */            -- # JMP
	/*     */            -- jmp_d:
	/* 110 */ 14x"2966", --     arg PC, GET_0
	/*     */            -- jmp_i:
	/* 111 */ 14x"0988", --     arg X, GET_0
	/* 112 */ 14x"0488", --     mem X, X, LOAD
	/* 113 */ 14x"2168", --     mov PC, X
	/*     */            -- jmp_cond_i:
	/* 114 */ 14x"0988", --     (-) arg X, GET_0
	/* 115 */ 14x"0488", --     (i) mem X, X, LOAD
	/* 116 */ 14x"3768", --     (-) cmv PC, X, COND_COPY
	/*     */            -- jmp_cond_d:
	/* 117 */ 14x"0988", --     (-) arg X, GET_0
	/* 118 */ 14x"3768", --     (-) cmv PC, X, COND_COPY
	/*     */            -- jmp_3dd:
	/* 119 */ 14x"0988", --     (--) arg X, GET_0
	/* 120 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 121 */ 14x"0baa", --     (--) arg Z, GET_2
	/* 122 */ 14x"1089", --     (--) cmp X, Y, UNSIGNED
	/* 123 */ 14x"376a", --     (--) cmv PC, Z, COND_COPY
	/*     */            -- jmp_3di:
	/* 124 */ 14x"0988", --     (--) arg X, GET_0
	/* 125 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 126 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 127 */ 14x"0baa", --     (--) arg Z, GET_2
	/* 128 */ 14x"1089", --     (--) cmp X, Y, UNSIGNED
	/* 129 */ 14x"376a", --     (--) cmv PC, Z, COND_COPY
	/*     */            -- jmp_3id:
	/* 130 */ 14x"0988", --     (--) arg X, GET_0
	/* 131 */ 14x"0488", --     (i-) mem X, X, LOAD
	/* 132 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 133 */ 14x"0baa", --     (--) arg Z, GET_2
	/* 134 */ 14x"1089", --     (--) cmp X, Y, UNSIGNED
	/* 135 */ 14x"376a", --     (--) cmv PC, Z, COND_COPY
	/*     */            -- jmp_3ii:
	/* 136 */ 14x"0988", --     (--) arg X, GET_0
	/* 137 */ 14x"0488", --     (i-) mem X, X, LOAD
	/* 138 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 139 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 140 */ 14x"0baa", --     (--) arg Z, GET_2
	/* 141 */ 14x"1089", --     (--) cmp X, Y, UNSIGNED
	/* 142 */ 14x"376a", --     (--) cmv PC, Z, COND_COPY
	/*     */            -- # ======================================
	/*     */            -- # MOV
	/*     */            -- mov_dd:
	/* 143 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 144 */ 14x"2899", --     (d-) arg Y, PUT
	/*     */            -- mov_di:
	/* 145 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 146 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 147 */ 14x"2899", --     (d-) arg Y, PUT
	/*     */            -- mov_id:
	/* 148 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 149 */ 14x"0988", --     (i-) arg X, GET_0
	/* 150 */ 14x"2589", --     (i-) mem X, Y, STORE
	/*     */            -- mov_ii:
	/* 151 */ 14x"0a99", --     (--) arg Y, GET_1
	/* 152 */ 14x"0499", --     (-i) mem Y, Y, LOAD
	/* 153 */ 14x"0988", --     (i-) arg X, GET_0
	/* 154 */ 14x"2589", --     (i-) mem X, Y, STORE
	/*     */            -- # ======================================
	/*     */            -- # Others
	/*     */            -- halt:
	/* 155 */ 14x"2166", --     mov PC, PC
	/*     */            -- getf:
	/* 156 */ 14x"2877", --     arg FL, PUT
	/*     */            -- setf:
	/* 157 */ 14x"0977", --     arg FL, GET_0
	/* 158 */ 14x"0284", --     con X, 0x3F # 6 bits
	/* 159 */ 14x"2e78", --     alu FL, X, AND
	/*     */            -- call_d:
	/* 160 */ 14x"0988", --     (-) arg X, GET_0
	/* 161 */ 14x"0d5c", --     (-) alu SP, 2, SUB
	/* 162 */ 14x"055d", --     (-) mem SP, NPC, STORE
	/* 163 */ 14x"2168", --     (-) mov PC, X
	/*     */            -- call_i:
	/* 164 */ 14x"0988", --     (-) arg X, GET_0
	/* 165 */ 14x"0488", --     (i) mem X, X, LOAD
	/* 166 */ 14x"0d5c", --     (-) alu SP, 2, SUB
	/* 167 */ 14x"055d", --     (-) mem SP, NPC, STORE
	/* 168 */ 14x"2168", --     (-) mov PC, X
	/*     */            -- ret:
	/* 169 */ 14x"0485", --     mem X, SP, LOAD
	/* 170 */ 14x"0c5c", --     alu SP, 2, ADD
	/* 171 */ 14x"2168", --     mov PC, X
	/*     */            -- push_d:
	/* 172 */ 14x"0988", --     (-) arg X, GET_0
	/* 173 */ 14x"0d5c", --     (-) alu SP, 2, SUB
	/* 174 */ 14x"2558", --     (-) mem SP, X, STORE
	/*     */            -- push_i:
	/* 175 */ 14x"0988", --     (-) arg X, GET_0
	/* 176 */ 14x"0488", --     (i) mem X, X, LOAD
	/* 177 */ 14x"0d5c", --     (-) alu SP, 2, SUB
	/* 178 */ 14x"2558", --     (-) mem SP, X, STORE
	/*     */            -- pop_d:
	/* 179 */ 14x"0495", --     (-) mem Y, SP, LOAD
	/* 180 */ 14x"0c5c", --     (-) alu SP, 2, ADD
	/* 181 */ 14x"2899", --     (d) arg Y, PUT
	/*     */            -- pop_i:
	/* 182 */ 14x"0495", --     (-) mem Y, SP, LOAD
	/* 183 */ 14x"0c5c", --     (-) alu SP, 2, ADD
	/* 184 */ 14x"0988", --     (i) arg X, GET_0
	/* 185 */ 14x"2589", --     (i) mem X, Y, STORE
	/*     */            -- mmap: # start, end, slot_idx / Y, Z, X
	/* 186 */ 14x"0999", --     arg, Y, GET_0
	/* 187 */ 14x"0aaa", --     arg, Z, GET_1
	/* 188 */ 14x"0b88", --     arg, X, GET_2
	/* 189 */ 14x"0300", --     mmu
	/* 190 */ 14x"01b6", --     mov K, PC
	/* 191 */ 14x"0160", --     mov PC, 0 # reset Fetcher
	/* 192 */ 14x"216b", --     mov PC, K
	/*     */            -- umap:
	/* 193 */ 14x"0988", --     arg, X, GET_0
	/* 194 */ 14x"0291", --     con Y, 0xFFFF
	/* 195 */ 14x"01a0", --     mov Z, 0
	/* 196 */ 14x"0300", --     mmu
	/* 197 */ 14x"01b6", --     mov K, PC
	/* 198 */ 14x"0160", --     mov PC, 0 # reset Fetcher
	/* 199 */ 14x"216b"  --     mov PC, K
	/*     */            -- end_of_uop_rom:
); -- uops_rom ---------------------------------------------------



constant label_reset : integer := 2;
constant label_alu_2dd : integer := 31;
constant label_alu_2di : integer := 35;
constant label_alu_2id : integer := 40;
constant label_alu_2ii : integer := 45;
constant label_alu_3dd : integer := 51;
constant label_alu_3di : integer := 55;
constant label_alu_3id : integer := 60;
constant label_alu_3ii : integer := 65;
constant label_alu_single_1dx : integer := 71;
constant label_alu_single_1ix : integer := 74;
constant label_alu_single_2dd : integer := 78;
constant label_alu_single_2di : integer := 81;
constant label_alu_single_2id : integer := 85;
constant label_alu_single_2ii : integer := 89;
constant label_cmp_dd : integer := 94;
constant label_cmp_di : integer := 97;
constant label_cmp_id : integer := 101;
constant label_cmp_ii : integer := 105;
constant label_jmp_d : integer := 110;
constant label_jmp_i : integer := 111;
constant label_jmp_cond_i : integer := 114;
constant label_jmp_cond_d : integer := 117;
constant label_jmp_3dd : integer := 119;
constant label_jmp_3di : integer := 124;
constant label_jmp_3id : integer := 130;
constant label_jmp_3ii : integer := 136;
constant label_mov_dd : integer := 143;
constant label_mov_di : integer := 145;
constant label_mov_id : integer := 148;
constant label_mov_ii : integer := 151;
constant label_halt : integer := 155;
constant label_getf : integer := 156;
constant label_setf : integer := 157;
constant label_call_d : integer := 160;
constant label_call_i : integer := 164;
constant label_ret : integer := 169;
constant label_push_d : integer := 172;
constant label_push_i : integer := 175;
constant label_pop_d : integer := 179;
constant label_pop_i : integer := 182;
constant label_mmap : integer := 186;
constant label_umap : integer := 193;
constant label_end_of_uop_rom : integer := 200;


type TArrUopsConstsROM is array (0 to 5-1) of TData;
constant uops_consts_rom : TArrUopsConstsROM := (
	x"0001", -- used 1 times
	x"FFFF", -- used 5 times
	x"00FF", -- used 1 times
	x"D000", -- used 2 times
	x"003F"  -- used 1 times
); -- uops_consts_rom -------------------------------------------

-- ##############################################################
-- ## END UOPS ROM
-- ##############################################################



