-- ##############################################################
-- ## BEGIN UOPS ROM
-- ##############################################################

type TArrUtopROM is array (0 to 25-1) of TUop;
signal uops_rom : TArrUtopROM := (
	"00000000000000", -- 0000 |     NULL # dummy instruction at index 0 & 1
	"00000000000000", -- 0000 |     NULL, FALLTHROUGH
	                  --      | reset:
	                  --      |     # reset arch registers
	"00000100010000", -- 0110 |     MOV A,  0
	"00000100100000", -- 0120 |     MOV B,  0
	"00000100110000", -- 0130 |     MOV C,  0
	"00000101000000", -- 0140 |     MOV D,  0
	"00000101010000", -- 0150 |     MOV SP, 0
	"00000101110000", -- 0170 |     MOV FL, 0
	"00000101100000", -- 0160 |     MOV PC, 0
	"00110101101101", -- 0d6d |     ALU PC, 2, SUB
	"00110101101101", -- 0d6d |     ALU PC, 2, SUB # reset vector PC=0xFFFB
	                  --      |     # reset MMU
	"00000110010000", -- 0190 |     MOV F, 0
	"00000110100000", -- 01a0 |     MOV G, 0
	"00110110101100", -- 0dac |     ALU G, 1, SUB
	"00000110000000", -- 0180 |     MOV E, 0
	"00001000000000", -- 0200 |     MMU # phy=A:B, idx=E, start=F, end=G
	"00000110100000", -- 01a0 |     MOV G, 0
	"00110010001100", -- 0c8c |     ALU E, 1, ADD
	"00001000000000", -- 0200 |     MMU # idx=1
	"00110010001100", -- 0c8c |     ALU E, 1, ADD
	"00001000000000", -- 0200 |     MMU # idx=2
	"00110010001100", -- 0c8c |     ALU E, 1, ADD
	"10001000000000", -- 2200 |     MMU # idx=3
	                  --      | alu2_ii:
	"10000100010000", -- 2110 |     MOV A,  0
	                  --      | alu2_ir:
	"10000100010000"  -- 2110 |     MOV A,  0
); -- uops_rom ---------------------------------------------------

constant uops_label_reset : integer := 2;
constant uops_label_alu2_ii : integer := 23;
constant uops_label_alu2_ir : integer := 24;

-- ##############################################################
-- ## END UOPS ROM
-- ##############################################################

